//
// Tangerine_top.v
//
// Top block for TangerineSDR Devkit version
// Start of block:  August 29, 2022
// Current version Date:
// Tom McDermott, N5EG
//

module Tangerine_top();

m10_rgmii eth0();

endmodule

